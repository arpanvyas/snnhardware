`include "header.vh"

module lookup_minus(
	input		clk,
	input		rst,
	input		[7:0]lut_in,
	output	[`W-1:0]lut_out
    );

wire		clk,rst;
wire		[7:0]lut_in;
reg		[`W-1:0]lut_out;


always @(posedge clk)
begin
	if (rst) begin
	lut_out =0;
	end else begin
	case (lut_in)
	
//		8'b00000001: lut_out = 24'b000000010010110000101100; //1
//		8'b00000010: lut_out = 24'b000000010110111010100001; //2
//		8'b00000011: lut_out = 24'b000000011011111111001101; //3
//		8'b00000100: lut_out = 24'b000000100010001011110010; //4
//		8'b00000101: lut_out = 24'b000000101001110000001011; //5
//		8'b00000110: lut_out = 24'b000000110010111111110011; //6
//		8'b00000111: lut_out = 24'b000000111110010010011011; //7
//		8'b00001000: lut_out = 24'b000001001100000101000001; //8
//		8'b00001001: lut_out = 24'b000001011100111011000010; //9
//		8'b00001010: lut_out = 24'b000001110001011111101111; //10
//		8'b00001011: lut_out = 24'b000010001010100111111100; //11
//		8'b00001100: lut_out = 24'b000010101001010100001110; //12
//		8'b00001101: lut_out = 24'b000011001110110011011001; //13
//		8'b00001110: lut_out = 24'b000011111100100101101111; //14
//		8'b00001111: lut_out = 24'b000100110100100000111000; //15
//		8'b00010000: lut_out = 24'b000101111000110100011101; //16
//		8'b00010001: lut_out = 24'b000111001100001111111010; //17
//		8'b00010010: lut_out = 24'b001000110010001001100001; //18
//		8'b00010011: lut_out = 24'b001010101110100111000011; //19
	

		8'b00010100: lut_out = 24'b000000000000000000001001; //-20
		8'b00010011: lut_out = 24'b000000000000000000001010; //-19
		8'b00010010: lut_out = 24'b000000000000000000001101; //-18
		8'b00010001: lut_out = 24'b000000000000000000010000; //-17
		8'b00010000: lut_out = 24'b000000000000000000010100; //-16
		8'b00001111: lut_out = 24'b000000000000000000011000; //-15
		8'b00001110: lut_out = 24'b000000000000000000011101; //-14
		8'b00001101: lut_out = 24'b000000000000000000100100; //-13
		8'b00001100: lut_out = 24'b000000000000000000101100; //-12
		8'b00001011: lut_out = 24'b000000000000000000110110; //-11
		8'b00001010: lut_out = 24'b000000000000000001000010; //-10
		8'b00001001: lut_out = 24'b000000000000000001010001; //-9
		8'b00001000: lut_out = 24'b000000000000000001100011; //-8
		8'b00000111: lut_out = 24'b000000000000000001111001; //-7
		8'b00000110: lut_out = 24'b000000000000000010010100; //-6
		8'b00000101: lut_out = 24'b000000000000000010110100; //-5
		8'b00000100: lut_out = 24'b000000000000000011011100; //-4
		8'b00000011: lut_out = 24'b000000000000000100001101; //-3
		8'b00000010: lut_out = 24'b000000000000000101001001; //-2	
	


		default	  : lut_out = 32'b000000000000000000000000;	
	endcase
	end
end 


//		8'b00010100: lut_out = 24'b000000000000000000001001; //-20
//		8'b00010011: lut_out = 24'b000000000000000000001010; //-19
//		8'b00010010: lut_out = 24'b000000000000000000001101; //-18
//		8'b00010001: lut_out = 24'b000000000000000000010000; //-17
//		8'b00010000: lut_out = 24'b000000000000000000010100; //-16
//		8'b00001111: lut_out = 24'b000000000000000000011000; //-15
//		8'b00001110: lut_out = 24'b000000000000000000011101; //-14
//		8'b00001101: lut_out = 24'b000000000000000000100100; //-13
//		8'b00001100: lut_out = 24'b000000000000000000101100; //-12
//		8'b00001011: lut_out = 24'b000000000000000000110110; //-11
//		8'b00001010: lut_out = 24'b000000000000000001000010; //-10
//		8'b00001001: lut_out = 24'b000000000000000001010001; //-9
//		8'b00001000: lut_out = 24'b000000000000000001100011; //-8
//		8'b00000111: lut_out = 24'b000000000000000001111001; //-7
//		8'b00000110: lut_out = 24'b000000000000000010010100; //-6
//		8'b00000101: lut_out = 24'b000000000000000010110100; //-5
//		8'b00000100: lut_out = 24'b000000000000000011011100; //-4
//		8'b00000011: lut_out = 24'b000000000000000100001101; //-3
//		8'b00000010: lut_out = 24'b000000000000000101001001; //-2



endmodule
