module rough(
    input clk,
    input  [9:0]ip,
    output [9:0] op
    );always@(posedge clk)
begin




end








endmodule
