`include "header.vh"

module lookup_plus(
	input		clk,
	input		rst,
	input		[7:0]lut_in,
	output	[23:0]lut_out
    );

wire		clk,rst;
wire		[7:0]lut_in;
reg		[23:0]lut_out;


always @(posedge clk)
begin
	if (rst) begin
	lut_out =0;
	end else begin
	case (lut_in)
	
//		8'b00010100: lut_out = 24'b111000001101000000010101; //-20
//		8'b00010011: lut_out = 24'b111001000111101000111000; //-19
//		8'b00010010: lut_out = 24'b111001111011011000011111; //-18
//		8'b00010001: lut_out = 24'b111010101001000010111101; //-17
//		8'b00010000: lut_out = 24'b111011010001010110000011; //-16
//		8'b00001111: lut_out = 24'b111011110100111010000101; //-15
//		8'b00001110: lut_out = 24'b111100010100010010101010; //-14
//		8'b00001101: lut_out = 24'b111100101111111111001111; //-13
//		8'b00001100: lut_out = 24'b111101001000011011100010; //-12
//		8'b00001011: lut_out = 24'b111101011110000000000001; //-11
//		8'b00001010: lut_out = 24'b111101110001000010010010; //-10
//		8'b00001001: lut_out = 24'b111110000001110101011010; //-9
//		8'b00001000: lut_out = 24'b111110010000101010001100; //-8
//		8'b00000111: lut_out = 24'b111110011101101111100000; //-7
//		8'b00000110: lut_out = 24'b111110101001010010011011; //-6
//		8'b00000101: lut_out = 24'b111110110011011110100001; //-5
//		8'b00000100: lut_out = 24'b111110111100011101111111; //-4
//		8'b00000011: lut_out = 24'b111111000100011001110101; //-3
//		8'b00000010: lut_out = 24'b111111001011011010000001; //-2
	
		8'b00000010: lut_out = 24'b111111111111111111101101; //2
		8'b00000011: lut_out = 24'b111111111111111111101010; //3
		8'b00000100: lut_out = 24'b111111111111111111100111; //4
		8'b00000101: lut_out = 24'b111111111111111111100100; //5
		8'b00000110: lut_out = 24'b111111111111111111100000; //6
		8'b00000111: lut_out = 24'b111111111111111111011100; //7
		8'b00001000: lut_out = 24'b111111111111111111010111; //8
		8'b00001001: lut_out = 24'b111111111111111111010010; //9
		8'b00001010: lut_out = 24'b111111111111111111001100; //10
		8'b00001011: lut_out = 24'b111111111111111111000101; //11
		8'b00001100: lut_out = 24'b111111111111111110111101; //12
		8'b00001101: lut_out = 24'b111111111111111110110100; //13
		8'b00001110: lut_out = 24'b111111111111111110101010; //14
		8'b00001111: lut_out = 24'b111111111111111110011111; //15
		8'b00010000: lut_out = 24'b111111111111111110010010; //16
		8'b00010001: lut_out = 24'b111111111111111110000011; //17
		8'b00010010: lut_out = 24'b111111111111111101110011; //18
		8'b00010011: lut_out = 24'b111111111111111101100000; //19
		8'b00010100: lut_out = 24'b111111111111111101001011; //20
//
//	8'b00010100: lut_out = 32'b11111110000011010000000101001011; //-20
//8'b00010011: lut_out = 32'b11111110010001111010001101110101; //-19
//8'b00010010: lut_out = 32'b11111110011110110110000111100010; //-18
//8'b00010001: lut_out = 32'b11111110101010010000101111001111; //-17
//8'b00010000: lut_out = 32'b11111110110100010101100000100010; //-16
//8'b00001111: lut_out = 32'b11111110111101001110100001000010; //-15
//8'b00001110: lut_out = 32'b11111111000101000100101010011111; //-14
//8'b00001101: lut_out = 32'b11111111001011111111110011101011; //-13
//8'b00001100: lut_out = 32'b11111111010010000110111000010110; //-12
//8'b00001011: lut_out = 32'b11111111010111100000000000000100; //-11
//8'b00001010: lut_out = 32'b11111111011100010000100100011010; //-10
//8'b00001001: lut_out = 32'b11111111100000011101010110010110; //-9
//8'b00001000: lut_out = 32'b11111111100100001010100011000000; //-8
//8'b00000111: lut_out = 32'b11111111100111011011110111111001; //-7
//8'b00000110: lut_out = 32'b11111111101010010100100110100110; //-6
//8'b00000101: lut_out = 32'b11111111101100110111101000000110; //-5
//8'b00000100: lut_out = 32'b11111111101111000111011111101000; //-4
//8'b00000011: lut_out = 32'b11111111110001000110011101010000; //-3
//8'b00000010: lut_out = 32'b11111111110010110110100000000101; //-2
	
	
	
	
//	
//8'b00010100: lut_out = 24'b110000011010000000101010; //-20
//8'b00010011: lut_out = 24'b110010001111010001110000; //-19
//8'b00010010: lut_out = 24'b110011110110110000111110; //-18
//8'b00010001: lut_out = 24'b110101010010000101111010; //-17
//8'b00010000: lut_out = 24'b110110100010101100000110; //-16
//8'b00001111: lut_out = 24'b110111101001110100001010; //-15
//8'b00001110: lut_out = 24'b111000101000100101010100; //-14
//8'b00001101: lut_out = 24'b111001011111111110011110; //-13
//8'b00001100: lut_out = 24'b111010010000110111000100; //-12
//8'b00001011: lut_out = 24'b111010111100000000000010; //-11
//8'b00001010: lut_out = 24'b111011100010000100100100; //-10
//8'b00001001: lut_out = 24'b111100000011101010110100; //-9
//8'b00001000: lut_out = 24'b111100100001010100011000; //-8
//8'b00000111: lut_out = 24'b111100111011011111000000; //-7
//8'b00000110: lut_out = 24'b111101010010100100110110; //-6
//8'b00000101: lut_out = 24'b111101100110111101000010; //-5
//8'b00000100: lut_out = 24'b111101111000111011111110; //-4
//8'b00000011: lut_out = 24'b111110001000110011101010; //-3
//8'b00000010: lut_out = 24'b111110010110110100000010; //-2


		default	  : lut_out = 24'b000000000000000000000000;	
	endcase
	end
end

//		8'b00000010: lut_out = 24'b111111111111111011010000; //2
//		8'b00000011: lut_out = 24'b111111111111111010100111; //3
//		8'b00000100: lut_out = 24'b111111111111111001111001; //4
//		8'b00000101: lut_out = 24'b111111111111111001000101; //5
//		8'b00000110: lut_out = 24'b111111111111111000001010; //6
//		8'b00000111: lut_out = 24'b111111111111110111000111; //7
//		8'b00001000: lut_out = 24'b111111111111110101111011; //8
//		8'b00001001: lut_out = 24'b111111111111110100100101; //9
//		8'b00001010: lut_out = 24'b111111111111110011000100; //10
//		8'b00001011: lut_out = 24'b111111111111110001010110; //11
//		8'b00001100: lut_out = 24'b111111111111101111011001; //12
//		8'b00001101: lut_out = 24'b111111111111101101001011; //13
//		8'b00001110: lut_out = 24'b111111111111101010101011; //14
//		8'b00001111: lut_out = 24'b111111111111100111110101; //15
//		8'b00010000: lut_out = 24'b111111111111100100100111; //16
//		8'b00010001: lut_out = 24'b111111111111100000111101; //17
//		8'b00010010: lut_out = 24'b111111111111011100110100; //18
//		8'b00010011: lut_out = 24'b111111111111011000001001; //19
//		8'b00010100: lut_out = 24'b111111111111010010110101; //20


endmodule
